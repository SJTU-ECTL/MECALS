module am8(input_A, input_B, product);
  wire [15:0] _000_;
  wire [15:0] _001_;
  wire [15:0] _002_;
  wire [15:0] _003_;
  wire [15:0] _004_;
  wire [15:0] _005_;
  wire [15:0] _006_;
  wire [15:0] _007_;
  wire [15:0] _008_;
  wire [15:0] _009_;
  wire [15:0] _010_;
  wire [15:0] _011_;
  wire [15:0] _012_;
  wire [15:0] _013_;
  wire [15:0] _014_;
  wire [15:0] _015_;
  wire [15:0] _016_;
  wire [15:0] _017_;
  wire [15:0] _018_;
  wire [15:0] _019_;
  wire [15:0] _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire [15:0] _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire [15:0] _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire [15:0] _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire [15:0] _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire [15:0] _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire [15:0] _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire [7:0] b0;
  wire [7:0] b1;
  wire [7:0] b2;
  wire [7:0] b3;
  wire [7:0] b4;
  wire [7:0] b5;
  wire [7:0] b6;
  wire [7:0] b7;
  input [7:0] input_A;
  input [7:0] input_B;
  wire [15:0] out;
  wire [7:0] pp1;
  wire [7:0] pp2;
  wire [7:0] pp3;
  wire [7:0] pp4;
  wire [7:0] pp5;
  wire [7:0] pp6;
  wire [7:0] pp7;
  wire [7:0] pp8;
  output [15:0] product;
  assign _001_[7] = _009_[7] ^ _008_[6];
  assign _001_[8] = _009_[8] ^ _008_[7];
  assign _001_[9] = _009_[9] ^ _008_[8];
  assign _001_[10] = _009_[10] ^ _008_[9];
  assign _001_[11] = _009_[11] ^ _008_[10];
  assign _001_[12] = _009_[12] ^ _008_[11];
  assign _001_[13] = _000_[13] ^ _008_[12];
  assign _001_[14] = _000_[14] ^ _008_[13];
  assign _001_[15] = _000_[15] ^ _008_[14];
  assign _001_[6] = pp7[0] ^ pp6[1];
  assign _009_[7] = _000_[7] ^ pp6[2];
  assign _009_[8] = _000_[8] ^ pp6[3];
  assign _009_[9] = _000_[9] ^ pp6[4];
  assign _009_[10] = _000_[10] ^ pp6[5];
  assign _009_[11] = _000_[11] ^ pp6[6];
  assign _009_[12] = _000_[12] ^ pp6[7];
  assign _008_[6] = pp7[0] & pp6[1];
  assign _039_[7] = _000_[7] & pp6[2];
  assign _039_[8] = _000_[8] & pp6[3];
  assign _039_[9] = _000_[9] & pp6[4];
  assign _039_[10] = _000_[10] & pp6[5];
  assign _039_[11] = _000_[11] & pp6[6];
  assign _039_[12] = _000_[12] & pp6[7];
  assign _002_[6] = _011_[6] ^ _010_[5];
  assign _002_[7] = _011_[7] ^ _010_[6];
  assign _002_[8] = _011_[8] ^ _010_[7];
  assign _002_[9] = _011_[9] ^ _010_[8];
  assign _002_[10] = _011_[10] ^ _010_[9];
  assign _002_[11] = _011_[11] ^ _010_[10];
  assign _002_[12] = _001_[12] ^ _010_[11];
  assign _002_[13] = _001_[13] ^ _010_[12];
  assign _002_[14] = _001_[14] ^ _010_[13];
  assign _002_[15] = _001_[15] ^ _010_[14];
  assign _002_[5] = pp6[0] ^ pp5[1];
  assign _011_[6] = _001_[6] ^ pp5[2];
  assign _011_[7] = _001_[7] ^ pp5[3];
  assign _011_[8] = _001_[8] ^ pp5[4];
  assign _011_[9] = _001_[9] ^ pp5[5];
  assign _011_[10] = _001_[10] ^ pp5[6];
  assign _011_[11] = _001_[11] ^ pp5[7];
  assign _010_[5] = pp6[0] & pp5[1];
  assign _058_[6] = _001_[6] & pp5[2];
  assign _058_[7] = _001_[7] & pp5[3];
  assign _058_[8] = _001_[8] & pp5[4];
  assign _058_[9] = _001_[9] & pp5[5];
  assign _058_[10] = _001_[10] & pp5[6];
  assign _058_[11] = _001_[11] & pp5[7];
  assign _003_[5] = _013_[5] ^ _012_[4];
  assign _003_[6] = _013_[6] ^ _012_[5];
  assign _003_[7] = _013_[7] ^ _012_[6];
  assign _003_[8] = _013_[8] ^ _012_[7];
  assign _003_[9] = _013_[9] ^ _012_[8];
  assign _003_[10] = _013_[10] ^ _012_[9];
  assign _003_[11] = _002_[11] ^ _012_[10];
  assign _003_[12] = _002_[12] ^ _012_[11];
  assign _003_[13] = _002_[13] ^ _012_[12];
  assign _003_[14] = _002_[14] ^ _012_[13];
  assign _003_[15] = _002_[15] ^ _012_[14];
  assign _003_[4] = pp5[0] ^ pp4[1];
  assign _013_[5] = _002_[5] ^ pp4[2];
  assign _013_[6] = _002_[6] ^ pp4[3];
  assign _013_[7] = _002_[7] ^ pp4[4];
  assign _013_[8] = _002_[8] ^ pp4[5];
  assign _013_[9] = _002_[9] ^ pp4[6];
  assign _013_[10] = _002_[10] ^ pp4[7];
  assign _012_[4] = pp5[0] & pp4[1];
  assign _078_[5] = _002_[5] & pp4[2];
  assign _078_[6] = _002_[6] & pp4[3];
  assign _078_[7] = _002_[7] & pp4[4];
  assign _078_[8] = _002_[8] & pp4[5];
  assign _078_[9] = _002_[9] & pp4[6];
  assign _078_[10] = _002_[10] & pp4[7];
  assign _004_[4] = _015_[4] ^ _014_[3];
  assign _004_[5] = _015_[5] ^ _014_[4];
  assign _004_[6] = _015_[6] ^ _014_[5];
  assign _004_[7] = _015_[7] ^ _014_[6];
  assign _004_[8] = _015_[8] ^ _014_[7];
  assign _004_[9] = _015_[9] ^ _014_[8];
  assign _004_[10] = _003_[10] ^ _014_[9];
  assign _004_[11] = _003_[11] ^ _014_[10];
  assign _004_[12] = _003_[12] ^ _014_[11];
  assign _004_[13] = _003_[13] ^ _014_[12];
  assign _004_[14] = _003_[14] ^ _014_[13];
  assign _004_[15] = _003_[15] ^ _014_[14];
  assign _004_[3] = pp4[0] ^ pp3[1];
  assign _015_[4] = _003_[4] ^ pp3[2];
  assign _015_[5] = _003_[5] ^ pp3[3];
  assign _015_[6] = _003_[6] ^ pp3[4];
  assign _015_[7] = _003_[7] ^ pp3[5];
  assign _015_[8] = _003_[8] ^ pp3[6];
  assign _015_[9] = _003_[9] ^ pp3[7];
  assign _014_[3] = pp4[0] & pp3[1];
  assign _098_[4] = _003_[4] & pp3[2];
  assign _098_[5] = _003_[5] & pp3[3];
  assign _098_[6] = _003_[6] & pp3[4];
  assign _098_[7] = _003_[7] & pp3[5];
  assign _098_[8] = _003_[8] & pp3[6];
  assign _098_[9] = _003_[9] & pp3[7];
  assign _005_[3] = _017_[3] ^ _016_[2];
  assign _005_[4] = _017_[4] ^ _016_[3];
  assign _005_[5] = _017_[5] ^ _016_[4];
  assign _005_[6] = _017_[6] ^ _016_[5];
  assign _005_[7] = _017_[7] ^ _016_[6];
  assign _005_[8] = _017_[8] ^ _016_[7];
  assign _005_[9] = _004_[9] ^ _016_[8];
  assign _005_[10] = _004_[10] ^ _016_[9];
  assign _005_[11] = _004_[11] ^ _016_[10];
  assign _005_[12] = _004_[12] ^ _016_[11];
  assign _005_[13] = _004_[13] ^ _016_[12];
  assign _005_[14] = _004_[14] ^ _016_[13];
  assign _005_[15] = _004_[15] ^ _016_[14];
  assign _005_[2] = pp3[0] ^ pp2[1];
  assign _017_[3] = _004_[3] ^ pp2[2];
  assign _017_[4] = _004_[4] ^ pp2[3];
  assign _017_[5] = _004_[5] ^ pp2[4];
  assign _017_[6] = _004_[6] ^ pp2[5];
  assign _017_[7] = _004_[7] ^ pp2[6];
  assign _017_[8] = _004_[8] ^ pp2[7];
  assign _016_[2] = pp3[0] & pp2[1];
  assign _122_[3] = _004_[3] & pp2[2];
  assign _122_[4] = _004_[4] & pp2[3];
  assign _122_[5] = _004_[5] & pp2[4];
  assign _122_[6] = _004_[6] & pp2[5];
  assign _122_[7] = _004_[7] & pp2[6];
  assign _122_[8] = _004_[8] & pp2[7];
  assign product[2] = _019_[2] ^ _018_[1];
  assign product[3] = _019_[3] ^ _018_[2];
  assign product[4] = _019_[4] ^ _018_[3];
  assign product[5] = _019_[5] ^ _018_[4];
  assign product[6] = _019_[6] ^ _018_[5];
  assign product[7] = _019_[7] ^ _018_[6];
  assign product[8] = _005_[8] ^ _018_[7];
  assign product[9] = _005_[9] ^ _018_[8];
  assign product[10] = _005_[10] ^ _018_[9];
  assign product[11] = _005_[11] ^ _018_[10];
  assign product[12] = _005_[12] ^ _018_[11];
  assign product[13] = _005_[13] ^ _018_[12];
  assign product[14] = _005_[14] ^ _018_[13];
  assign product[15] = _005_[15] ^ _018_[14];
  assign product[1] = pp1[1] ^ pp2[0];
  assign _019_[2] = pp1[2] ^ _005_[2];
  assign _019_[3] = pp1[3] ^ _005_[3];
  assign _019_[4] = pp1[4] ^ _005_[4];
  assign _019_[5] = pp1[5] ^ _005_[5];
  assign _019_[6] = pp1[6] ^ _005_[6];
  assign _019_[7] = pp1[7] ^ _005_[7];
  assign _018_[1] = pp1[1] & pp2[0];
  assign _146_[2] = pp1[2] & _005_[2];
  assign _146_[3] = pp1[3] & _005_[3];
  assign _146_[4] = pp1[4] & _005_[4];
  assign _146_[5] = pp1[5] & _005_[5];
  assign _146_[6] = pp1[6] & _005_[6];
  assign _146_[7] = pp1[7] & _005_[7];
  assign pp2[0] = input_A[0] & input_B[1];
  assign pp2[1] = input_A[1] & input_B[1];
  assign pp2[2] = input_A[2] & input_B[1];
  assign pp2[3] = input_A[3] & input_B[1];
  assign pp2[4] = input_A[4] & input_B[1];
  assign pp2[5] = input_A[5] & input_B[1];
  assign pp2[6] = input_A[6] & input_B[1];
  assign pp2[7] = input_A[7] & input_B[1];
  assign _021_ = _007_[9] & _020_[8];
  assign _022_ = _007_[11] & _020_[10];
  assign _023_ = _007_[13] & _020_[12];
  assign pp3[0] = input_A[0] & input_B[2];
  assign _024_ = _026_ & _035_;
  assign pp3[1] = input_A[1] & input_B[2];
  assign _025_ = _007_[9] & _007_[8];
  assign _026_ = _007_[11] & _007_[10];
  assign _027_ = _007_[13] & _007_[12];
  assign _028_ = _026_ & _025_;
  assign pp3[2] = input_A[2] & input_B[2];
  assign _029_ = _028_ & _006_[7];
  assign _030_ = _025_ & _006_[7];
  assign _031_ = _027_ & _006_[11];
  assign pp3[3] = input_A[3] & input_B[2];
  assign _032_ = _007_[8] & _006_[7];
  assign _033_ = _007_[10] & _006_[9];
  assign _034_ = _007_[12] & _006_[11];
  assign _000_[15] = pp8[7] & _006_[13];
  assign _035_ = _020_[9] | _021_;
  assign _036_ = _020_[11] | _022_;
  assign _037_ = _020_[13] | _023_;
  assign pp3[4] = input_A[4] & input_B[2];
  assign _038_ = _036_ | _024_;
  assign pp3[5] = input_A[5] & input_B[2];
  assign _006_[11] = _038_ | _029_;
  assign _006_[9] = _035_ | _030_;
  assign _006_[13] = _037_ | _031_;
  assign _006_[8] = _020_[8] | _032_;
  assign _006_[10] = _020_[10] | _033_;
  assign _006_[12] = _020_[12] | _034_;
  assign pp3[6] = input_A[6] & input_B[2];
  assign _040_ = _009_[9] & _039_[8];
  assign _041_ = _009_[11] & _039_[10];
  assign _042_ = _000_[13] & _039_[12];
  assign _043_ = _046_ & _055_;
  assign pp3[7] = input_A[7] & input_B[2];
  assign _044_ = _009_[7] & _008_[6];
  assign _045_ = _009_[9] & _009_[8];
  assign _046_ = _009_[11] & _009_[10];
  assign pp4[0] = input_A[0] & input_B[3];
  assign _047_ = _000_[13] & _009_[12];
  assign _048_ = _046_ & _045_;
  assign _049_ = _048_ & _008_[7];
  assign pp4[1] = input_A[1] & input_B[3];
  assign _050_ = _045_ & _008_[7];
  assign _051_ = _047_ & _008_[11];
  assign _052_ = _009_[8] & _008_[7];
  assign _053_ = _009_[10] & _008_[9];
  assign _054_ = _009_[12] & _008_[11];
  assign _008_[14] = _000_[14] & _008_[13];
  assign pp4[2] = input_A[2] & input_B[3];
  assign _055_ = _039_[9] | _040_;
  assign _056_ = _039_[11] | _041_;
  assign _057_ = _056_ | _043_;
  assign pp4[3] = input_A[3] & input_B[3];
  assign _008_[7] = _039_[7] | _044_;
  assign _008_[11] = _057_ | _049_;
  assign _008_[9] = _055_ | _050_;
  assign _008_[13] = _042_ | _051_;
  assign pp4[4] = input_A[4] & input_B[3];
  assign _008_[8] = _039_[8] | _052_;
  assign _008_[10] = _039_[10] | _053_;
  assign _008_[12] = _039_[12] | _054_;
  assign _059_ = _011_[9] & _058_[8];
  assign _060_ = _011_[11] & _058_[10];
  assign pp4[5] = input_A[5] & input_B[3];
  assign _061_ = _064_ & _010_[5];
  assign _062_ = _066_ & _074_;
  assign pp4[6] = input_A[6] & input_B[3];
  assign _063_ = _011_[7] & _058_[6];
  assign _064_ = _011_[7] & _011_[6];
  assign _065_ = _011_[9] & _011_[8];
  assign _066_ = _011_[11] & _011_[10];
  assign _067_ = _001_[13] & _001_[12];
  assign _068_ = _066_ & _065_;
  assign pp4[7] = input_A[7] & input_B[3];
  assign _069_ = _068_ & _010_[7];
  assign _070_ = _065_ & _010_[7];
  assign _010_[13] = _067_ & _010_[11];
  assign _071_ = _011_[6] & _010_[5];
  assign pp5[0] = input_A[0] & input_B[4];
  assign _072_ = _011_[8] & _010_[7];
  assign _073_ = _011_[10] & _010_[9];
  assign _010_[12] = _001_[12] & _010_[11];
  assign _010_[14] = _001_[14] & _010_[13];
  assign _074_ = _058_[9] | _059_;
  assign _075_ = _058_[11] | _060_;
  assign pp5[1] = input_A[1] & input_B[4];
  assign _010_[7] = _077_ | _061_;
  assign _076_ = _075_ | _062_;
  assign _077_ = _058_[7] | _063_;
  assign pp5[2] = input_A[2] & input_B[4];
  assign _010_[11] = _076_ | _069_;
  assign _010_[9] = _074_ | _070_;
  assign _010_[6] = _058_[6] | _071_;
  assign _010_[8] = _058_[8] | _072_;
  assign _010_[10] = _058_[10] | _073_;
  assign pp5[3] = input_A[3] & input_B[4];
  assign _079_ = _013_[9] & _078_[8];
  assign _080_ = _002_[11] & _078_[10];
  assign _081_ = _085_ & _012_[5];
  assign _082_ = _087_ & _095_;
  assign pp5[4] = input_A[4] & input_B[4];
  assign _083_ = _013_[5] & _012_[4];
  assign _084_ = _013_[7] & _078_[6];
  assign _085_ = _013_[7] & _013_[6];
  assign _086_ = _013_[9] & _013_[8];
  assign _087_ = _002_[11] & _013_[10];
  assign pp5[5] = input_A[5] & input_B[4];
  assign _088_ = _002_[13] & _002_[12];
  assign _089_ = _087_ & _086_;
  assign _090_ = _089_ & _012_[7];
  assign pp5[6] = input_A[6] & input_B[4];
  assign _091_ = _086_ & _012_[7];
  assign _012_[13] = _088_ & _012_[11];
  assign _092_ = _013_[6] & _012_[5];
  assign _093_ = _013_[8] & _012_[7];
  assign _094_ = _013_[10] & _012_[9];
  assign _012_[12] = _002_[12] & _012_[11];
  assign _012_[14] = _002_[14] & _012_[13];
  assign pp5[7] = input_A[7] & input_B[4];
  assign _095_ = _078_[9] | _079_;
  assign _012_[7] = _097_ | _081_;
  assign _096_ = _080_ | _082_;
  assign pp6[0] = input_A[0] & input_B[5];
  assign _012_[5] = _078_[5] | _083_;
  assign _097_ = _078_[7] | _084_;
  assign _012_[11] = _096_ | _090_;
  assign _012_[9] = _095_ | _091_;
  assign pp6[1] = input_A[1] & input_B[5];
  assign _012_[6] = _078_[6] | _092_;
  assign _012_[8] = _078_[8] | _093_;
  assign _012_[10] = _078_[10] | _094_;
  assign _099_ = _015_[9] & _098_[8];
  assign pp6[2] = input_A[2] & input_B[5];
  assign _100_ = _105_ & _120_;
  assign _101_ = _107_ & _118_;
  assign _102_ = _109_ & _014_[3];
  assign pp6[3] = input_A[3] & input_B[5];
  assign _103_ = _015_[5] & _098_[4];
  assign _104_ = _015_[7] & _098_[6];
  assign _105_ = _015_[7] & _015_[6];
  assign _106_ = _015_[9] & _015_[8];
  assign _107_ = _003_[11] & _003_[10];
  assign _108_ = _003_[13] & _003_[12];
  assign _109_ = _105_ & _111_;
  assign _110_ = _107_ & _106_;
  assign pp6[4] = input_A[4] & input_B[5];
  assign _111_ = _015_[5] & _015_[4];
  assign _112_ = _110_ & _014_[7];
  assign _113_ = _111_ & _014_[3];
  assign _114_ = _106_ & _014_[7];
  assign _014_[13] = _108_ & _014_[11];
  assign _115_ = _015_[4] & _014_[3];
  assign _116_ = _015_[6] & _014_[5];
  assign pp6[5] = input_A[5] & input_B[5];
  assign _117_ = _015_[8] & _014_[7];
  assign _014_[10] = _003_[10] & _014_[9];
  assign _014_[12] = _003_[12] & _014_[11];
  assign _014_[14] = _003_[14] & _014_[13];
  assign _118_ = _098_[9] | _099_;
  assign pp6[6] = input_A[6] & input_B[5];
  assign _119_ = _121_ | _100_;
  assign _014_[7] = _119_ | _102_;
  assign _120_ = _098_[5] | _103_;
  assign _121_ = _098_[7] | _104_;
  assign pp6[7] = input_A[7] & input_B[5];
  assign _014_[11] = _101_ | _112_;
  assign _014_[5] = _120_ | _113_;
  assign _014_[9] = _118_ | _114_;
  assign _014_[4] = _098_[4] | _115_;
  assign _014_[6] = _098_[6] | _116_;
  assign _014_[8] = _098_[8] | _117_;
  assign pp7[0] = input_A[0] & input_B[6];
  assign _123_ = _004_[9] & _122_[8];
  assign _124_ = _130_ & _144_;
  assign _125_ = _132_ & _123_;
  assign pp7[1] = input_A[1] & input_B[6];
  assign _126_ = _134_ & _016_[3];
  assign _127_ = _017_[3] & _016_[2];
  assign _128_ = _017_[5] & _122_[4];
  assign _129_ = _017_[7] & _122_[6];
  assign _130_ = _017_[7] & _017_[6];
  assign _131_ = _004_[9] & _017_[8];
  assign _132_ = _004_[11] & _004_[10];
  assign pp7[2] = input_A[2] & input_B[6];
  assign _133_ = _004_[13] & _004_[12];
  assign _134_ = _130_ & _136_;
  assign _135_ = _132_ & _131_;
  assign _136_ = _017_[5] & _017_[4];
  assign _137_ = _135_ & _016_[7];
  assign _138_ = _136_ & _016_[3];
  assign pp7[3] = input_A[3] & input_B[6];
  assign _139_ = _131_ & _016_[7];
  assign _016_[13] = _133_ & _016_[11];
  assign _140_ = _017_[4] & _016_[3];
  assign _141_ = _017_[6] & _016_[5];
  assign _142_ = _017_[8] & _016_[7];
  assign _016_[10] = _004_[10] & _016_[9];
  assign _016_[12] = _004_[12] & _016_[11];
  assign _016_[14] = _004_[14] & _016_[13];
  assign pp7[4] = input_A[4] & input_B[6];
  assign _143_ = _145_ | _124_;
  assign _016_[7] = _143_ | _126_;
  assign pp7[5] = input_A[5] & input_B[6];
  assign _016_[3] = _122_[3] | _127_;
  assign _144_ = _122_[5] | _128_;
  assign _145_ = _122_[7] | _129_;
  assign _016_[11] = _125_ | _137_;
  assign _016_[5] = _144_ | _138_;
  assign _016_[9] = _123_ | _139_;
  assign pp7[6] = input_A[6] & input_B[6];
  assign _016_[4] = _122_[4] | _140_;
  assign _016_[6] = _122_[6] | _141_;
  assign _016_[8] = _122_[8] | _142_;
  assign pp7[7] = input_A[7] & input_B[6];
  assign _147_ = _159_ & _018_[1];
  assign _148_ = _153_ & _167_;
  assign _149_ = _157_ & _018_[3];
  assign _150_ = _019_[3] & _146_[2];
  assign pp8[0] = input_A[0] & input_B[7];
  assign _151_ = _019_[5] & _146_[4];
  assign _152_ = _019_[7] & _146_[6];
  assign _153_ = _019_[7] & _019_[6];
  assign _154_ = _005_[9] & _005_[8];
  assign _155_ = _005_[11] & _005_[10];
  assign _156_ = _005_[13] & _005_[12];
  assign _157_ = _153_ & _160_;
  assign _158_ = _155_ & _154_;
  assign pp8[1] = input_A[1] & input_B[7];
  assign _159_ = _019_[3] & _019_[2];
  assign _160_ = _019_[5] & _019_[4];
  assign _018_[11] = _158_ & _018_[7];
  assign _161_ = _160_ & _018_[3];
  assign _018_[9] = _154_ & _018_[7];
  assign _018_[13] = _156_ & _018_[11];
  assign _162_ = _019_[2] & _018_[1];
  assign _163_ = _019_[4] & _018_[3];
  assign _164_ = _019_[6] & _018_[5];
  assign pp8[2] = input_A[2] & input_B[7];
  assign _018_[8] = _005_[8] & _018_[7];
  assign _018_[10] = _005_[10] & _018_[9];
  assign _018_[12] = _005_[12] & _018_[11];
  assign _018_[14] = _005_[14] & _018_[13];
  assign _018_[3] = _166_ | _147_;
  assign pp8[3] = input_A[3] & input_B[7];
  assign _165_ = _168_ | _148_;
  assign _018_[7] = _165_ | _149_;
  assign _166_ = _146_[3] | _150_;
  assign _167_ = _146_[5] | _151_;
  assign _168_ = _146_[7] | _152_;
  assign pp8[4] = input_A[4] & input_B[7];
  assign _018_[5] = _167_ | _161_;
  assign _018_[2] = _146_[2] | _162_;
  assign _018_[4] = _146_[4] | _163_;
  assign _018_[6] = _146_[6] | _164_;
  assign pp8[5] = input_A[5] & input_B[7];
  assign pp8[6] = input_A[6] & input_B[7];
  assign pp8[7] = input_A[7] & input_B[7];
  assign product[0] = input_A[0] & input_B[0];
  assign pp1[1] = input_A[1] & input_B[0];
  assign pp1[2] = input_A[2] & input_B[0];
  assign pp1[3] = input_A[3] & input_B[0];
  assign pp1[4] = input_A[4] & input_B[0];
  assign pp1[5] = input_A[5] & input_B[0];
  assign pp1[6] = input_A[6] & input_B[0];
  assign pp1[7] = input_A[7] & input_B[0];
  assign _000_[8] = _007_[8] ^ _006_[7];
  assign _000_[9] = _007_[9] ^ _006_[8];
  assign _000_[10] = _007_[10] ^ _006_[9];
  assign _000_[11] = _007_[11] ^ _006_[10];
  assign _000_[12] = _007_[12] ^ _006_[11];
  assign _000_[13] = _007_[13] ^ _006_[12];
  assign _000_[14] = pp8[7] ^ _006_[13];
  assign _000_[7] = pp8[0] ^ pp7[1];
  assign _007_[8] = pp8[1] ^ pp7[2];
  assign _007_[9] = pp8[2] ^ pp7[3];
  assign _007_[10] = pp8[3] ^ pp7[4];
  assign _007_[11] = pp8[4] ^ pp7[5];
  assign _007_[12] = pp8[5] ^ pp7[6];
  assign _007_[13] = pp8[6] ^ pp7[7];
  assign _006_[7] = pp8[0] & pp7[1];
  assign _020_[8] = pp8[1] & pp7[2];
  assign _020_[9] = pp8[2] & pp7[3];
  assign _020_[10] = pp8[3] & pp7[4];
  assign _020_[11] = pp8[4] & pp7[5];
  assign _020_[12] = pp8[5] & pp7[6];
  assign _020_[13] = pp8[6] & pp7[7];
  assign _000_[6:0] = { pp7[0], 6'h00 };
  assign _001_[5:0] = { pp6[0], 5'h00 };
  assign _002_[4:0] = { pp5[0], 4'h0 };
  assign _003_[3:0] = { pp4[0], 3'h0 };
  assign _004_[2:0] = { pp3[0], 2'h0 };
  assign _005_[1:0] = { pp2[0], 1'h0 };
  assign { _006_[15:14], _006_[6:0] } = { 1'h0, _000_[15], 7'h00 };
  assign { _007_[15:14], _007_[7:0] } = { 1'h0, pp8[7], _000_[7], pp7[0], 6'h00 };
  assign _008_[5:0] = 6'h00;
  assign { _009_[15:13], _009_[6:0] } = { _000_[15:13], _001_[6], pp6[0], 5'h00 };
  assign _010_[4:0] = 5'h00;
  assign { _011_[15:12], _011_[5:0] } = { _001_[15:12], _002_[5], pp5[0], 4'h0 };
  assign _012_[3:0] = 4'h0;
  assign { _013_[15:11], _013_[4:0] } = { _002_[15:11], _003_[4], pp4[0], 3'h0 };
  assign _014_[2:0] = 3'h0;
  assign { _015_[15:10], _015_[3:0] } = { _003_[15:10], _004_[3], pp3[0], 2'h0 };
  assign _016_[1:0] = 2'h0;
  assign { _017_[15:9], _017_[2:0] } = { _004_[15:9], _005_[2], pp2[0], 1'h0 };
  assign _018_[0] = 1'h0;
  assign { _019_[15:8], _019_[1:0] } = { _005_[15:8], product[1:0] };
  assign { _020_[15:14], _020_[7:0] } = { 2'h0, _006_[7], 7'h00 };
  assign { _039_[15:13], _039_[6:0] } = { 3'h0, _008_[6], 6'h00 };
  assign { _058_[15:12], _058_[5:0] } = { 4'h0, _010_[5], 5'h00 };
  assign { _078_[15:11], _078_[4:0] } = { 5'h00, _012_[4], 4'h0 };
  assign { _098_[15:10], _098_[3:0] } = { 6'h00, _014_[3], 3'h0 };
  assign { _122_[15:9], _122_[2:0] } = { 7'h00, _016_[2], 2'h0 };
  assign { _146_[15:8], _146_[1:0] } = { 8'h00, _018_[1], 1'h0 };
  assign b0 = { 7'h00, input_B[0] };
  assign b1 = { 7'h00, input_B[1] };
  assign b2 = { 7'h00, input_B[2] };
  assign b3 = { 7'h00, input_B[3] };
  assign b4 = { 7'h00, input_B[4] };
  assign b5 = { 7'h00, input_B[5] };
  assign b6 = { 7'h00, input_B[6] };
  assign b7 = { 7'h00, input_B[7] };
  assign out = product;
  assign pp1[0] = product[0];
endmodule
