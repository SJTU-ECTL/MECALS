module rca32(input_A, input_B, output_sum);
  wire \adder[0].adder_inst.in_A ;
  wire \adder[0].adder_inst.in_B ;
  wire \adder[0].adder_inst.in_carry ;
  wire \adder[0].adder_inst.intermediateResult1 ;
  wire \adder[0].adder_inst.intermediateResult2 ;
  wire \adder[0].adder_inst.intermediateResult3 ;
  wire \adder[0].adder_inst.out_carry ;
  wire \adder[0].adder_inst.out_sum ;
  wire \adder[10].adder_inst.in_A ;
  wire \adder[10].adder_inst.in_B ;
  wire \adder[10].adder_inst.in_carry ;
  wire \adder[10].adder_inst.intermediateResult1 ;
  wire \adder[10].adder_inst.intermediateResult2 ;
  wire \adder[10].adder_inst.intermediateResult3 ;
  wire \adder[10].adder_inst.out_carry ;
  wire \adder[10].adder_inst.out_sum ;
  wire \adder[11].adder_inst.in_A ;
  wire \adder[11].adder_inst.in_B ;
  wire \adder[11].adder_inst.in_carry ;
  wire \adder[11].adder_inst.intermediateResult1 ;
  wire \adder[11].adder_inst.intermediateResult2 ;
  wire \adder[11].adder_inst.intermediateResult3 ;
  wire \adder[11].adder_inst.out_carry ;
  wire \adder[11].adder_inst.out_sum ;
  wire \adder[12].adder_inst.in_A ;
  wire \adder[12].adder_inst.in_B ;
  wire \adder[12].adder_inst.in_carry ;
  wire \adder[12].adder_inst.intermediateResult1 ;
  wire \adder[12].adder_inst.intermediateResult2 ;
  wire \adder[12].adder_inst.intermediateResult3 ;
  wire \adder[12].adder_inst.out_carry ;
  wire \adder[12].adder_inst.out_sum ;
  wire \adder[13].adder_inst.in_A ;
  wire \adder[13].adder_inst.in_B ;
  wire \adder[13].adder_inst.in_carry ;
  wire \adder[13].adder_inst.intermediateResult1 ;
  wire \adder[13].adder_inst.intermediateResult2 ;
  wire \adder[13].adder_inst.intermediateResult3 ;
  wire \adder[13].adder_inst.out_carry ;
  wire \adder[13].adder_inst.out_sum ;
  wire \adder[14].adder_inst.in_A ;
  wire \adder[14].adder_inst.in_B ;
  wire \adder[14].adder_inst.in_carry ;
  wire \adder[14].adder_inst.intermediateResult1 ;
  wire \adder[14].adder_inst.intermediateResult2 ;
  wire \adder[14].adder_inst.intermediateResult3 ;
  wire \adder[14].adder_inst.out_carry ;
  wire \adder[14].adder_inst.out_sum ;
  wire \adder[15].adder_inst.in_A ;
  wire \adder[15].adder_inst.in_B ;
  wire \adder[15].adder_inst.in_carry ;
  wire \adder[15].adder_inst.intermediateResult1 ;
  wire \adder[15].adder_inst.intermediateResult2 ;
  wire \adder[15].adder_inst.intermediateResult3 ;
  wire \adder[15].adder_inst.out_carry ;
  wire \adder[15].adder_inst.out_sum ;
  wire \adder[16].adder_inst.in_A ;
  wire \adder[16].adder_inst.in_B ;
  wire \adder[16].adder_inst.in_carry ;
  wire \adder[16].adder_inst.intermediateResult1 ;
  wire \adder[16].adder_inst.intermediateResult2 ;
  wire \adder[16].adder_inst.intermediateResult3 ;
  wire \adder[16].adder_inst.out_carry ;
  wire \adder[16].adder_inst.out_sum ;
  wire \adder[17].adder_inst.in_A ;
  wire \adder[17].adder_inst.in_B ;
  wire \adder[17].adder_inst.in_carry ;
  wire \adder[17].adder_inst.intermediateResult1 ;
  wire \adder[17].adder_inst.intermediateResult2 ;
  wire \adder[17].adder_inst.intermediateResult3 ;
  wire \adder[17].adder_inst.out_carry ;
  wire \adder[17].adder_inst.out_sum ;
  wire \adder[18].adder_inst.in_A ;
  wire \adder[18].adder_inst.in_B ;
  wire \adder[18].adder_inst.in_carry ;
  wire \adder[18].adder_inst.intermediateResult1 ;
  wire \adder[18].adder_inst.intermediateResult2 ;
  wire \adder[18].adder_inst.intermediateResult3 ;
  wire \adder[18].adder_inst.out_carry ;
  wire \adder[18].adder_inst.out_sum ;
  wire \adder[19].adder_inst.in_A ;
  wire \adder[19].adder_inst.in_B ;
  wire \adder[19].adder_inst.in_carry ;
  wire \adder[19].adder_inst.intermediateResult1 ;
  wire \adder[19].adder_inst.intermediateResult2 ;
  wire \adder[19].adder_inst.intermediateResult3 ;
  wire \adder[19].adder_inst.out_carry ;
  wire \adder[19].adder_inst.out_sum ;
  wire \adder[1].adder_inst.in_A ;
  wire \adder[1].adder_inst.in_B ;
  wire \adder[1].adder_inst.in_carry ;
  wire \adder[1].adder_inst.intermediateResult1 ;
  wire \adder[1].adder_inst.intermediateResult2 ;
  wire \adder[1].adder_inst.intermediateResult3 ;
  wire \adder[1].adder_inst.out_carry ;
  wire \adder[1].adder_inst.out_sum ;
  wire \adder[20].adder_inst.in_A ;
  wire \adder[20].adder_inst.in_B ;
  wire \adder[20].adder_inst.in_carry ;
  wire \adder[20].adder_inst.intermediateResult1 ;
  wire \adder[20].adder_inst.intermediateResult2 ;
  wire \adder[20].adder_inst.intermediateResult3 ;
  wire \adder[20].adder_inst.out_carry ;
  wire \adder[20].adder_inst.out_sum ;
  wire \adder[21].adder_inst.in_A ;
  wire \adder[21].adder_inst.in_B ;
  wire \adder[21].adder_inst.in_carry ;
  wire \adder[21].adder_inst.intermediateResult1 ;
  wire \adder[21].adder_inst.intermediateResult2 ;
  wire \adder[21].adder_inst.intermediateResult3 ;
  wire \adder[21].adder_inst.out_carry ;
  wire \adder[21].adder_inst.out_sum ;
  wire \adder[22].adder_inst.in_A ;
  wire \adder[22].adder_inst.in_B ;
  wire \adder[22].adder_inst.in_carry ;
  wire \adder[22].adder_inst.intermediateResult1 ;
  wire \adder[22].adder_inst.intermediateResult2 ;
  wire \adder[22].adder_inst.intermediateResult3 ;
  wire \adder[22].adder_inst.out_carry ;
  wire \adder[22].adder_inst.out_sum ;
  wire \adder[23].adder_inst.in_A ;
  wire \adder[23].adder_inst.in_B ;
  wire \adder[23].adder_inst.in_carry ;
  wire \adder[23].adder_inst.intermediateResult1 ;
  wire \adder[23].adder_inst.intermediateResult2 ;
  wire \adder[23].adder_inst.intermediateResult3 ;
  wire \adder[23].adder_inst.out_carry ;
  wire \adder[23].adder_inst.out_sum ;
  wire \adder[24].adder_inst.in_A ;
  wire \adder[24].adder_inst.in_B ;
  wire \adder[24].adder_inst.in_carry ;
  wire \adder[24].adder_inst.intermediateResult1 ;
  wire \adder[24].adder_inst.intermediateResult2 ;
  wire \adder[24].adder_inst.intermediateResult3 ;
  wire \adder[24].adder_inst.out_carry ;
  wire \adder[24].adder_inst.out_sum ;
  wire \adder[25].adder_inst.in_A ;
  wire \adder[25].adder_inst.in_B ;
  wire \adder[25].adder_inst.in_carry ;
  wire \adder[25].adder_inst.intermediateResult1 ;
  wire \adder[25].adder_inst.intermediateResult2 ;
  wire \adder[25].adder_inst.intermediateResult3 ;
  wire \adder[25].adder_inst.out_carry ;
  wire \adder[25].adder_inst.out_sum ;
  wire \adder[26].adder_inst.in_A ;
  wire \adder[26].adder_inst.in_B ;
  wire \adder[26].adder_inst.in_carry ;
  wire \adder[26].adder_inst.intermediateResult1 ;
  wire \adder[26].adder_inst.intermediateResult2 ;
  wire \adder[26].adder_inst.intermediateResult3 ;
  wire \adder[26].adder_inst.out_carry ;
  wire \adder[26].adder_inst.out_sum ;
  wire \adder[27].adder_inst.in_A ;
  wire \adder[27].adder_inst.in_B ;
  wire \adder[27].adder_inst.in_carry ;
  wire \adder[27].adder_inst.intermediateResult1 ;
  wire \adder[27].adder_inst.intermediateResult2 ;
  wire \adder[27].adder_inst.intermediateResult3 ;
  wire \adder[27].adder_inst.out_carry ;
  wire \adder[27].adder_inst.out_sum ;
  wire \adder[28].adder_inst.in_A ;
  wire \adder[28].adder_inst.in_B ;
  wire \adder[28].adder_inst.in_carry ;
  wire \adder[28].adder_inst.intermediateResult1 ;
  wire \adder[28].adder_inst.intermediateResult2 ;
  wire \adder[28].adder_inst.intermediateResult3 ;
  wire \adder[28].adder_inst.out_carry ;
  wire \adder[28].adder_inst.out_sum ;
  wire \adder[29].adder_inst.in_A ;
  wire \adder[29].adder_inst.in_B ;
  wire \adder[29].adder_inst.in_carry ;
  wire \adder[29].adder_inst.intermediateResult1 ;
  wire \adder[29].adder_inst.intermediateResult2 ;
  wire \adder[29].adder_inst.intermediateResult3 ;
  wire \adder[29].adder_inst.out_carry ;
  wire \adder[29].adder_inst.out_sum ;
  wire \adder[2].adder_inst.in_A ;
  wire \adder[2].adder_inst.in_B ;
  wire \adder[2].adder_inst.in_carry ;
  wire \adder[2].adder_inst.intermediateResult1 ;
  wire \adder[2].adder_inst.intermediateResult2 ;
  wire \adder[2].adder_inst.intermediateResult3 ;
  wire \adder[2].adder_inst.out_carry ;
  wire \adder[2].adder_inst.out_sum ;
  wire \adder[30].adder_inst.in_A ;
  wire \adder[30].adder_inst.in_B ;
  wire \adder[30].adder_inst.in_carry ;
  wire \adder[30].adder_inst.intermediateResult1 ;
  wire \adder[30].adder_inst.intermediateResult2 ;
  wire \adder[30].adder_inst.intermediateResult3 ;
  wire \adder[30].adder_inst.out_carry ;
  wire \adder[30].adder_inst.out_sum ;
  wire \adder[31].adder_inst.in_A ;
  wire \adder[31].adder_inst.in_B ;
  wire \adder[31].adder_inst.in_carry ;
  wire \adder[31].adder_inst.intermediateResult1 ;
  wire \adder[31].adder_inst.intermediateResult2 ;
  wire \adder[31].adder_inst.intermediateResult3 ;
  wire \adder[31].adder_inst.out_carry ;
  wire \adder[31].adder_inst.out_sum ;
  wire \adder[3].adder_inst.in_A ;
  wire \adder[3].adder_inst.in_B ;
  wire \adder[3].adder_inst.in_carry ;
  wire \adder[3].adder_inst.intermediateResult1 ;
  wire \adder[3].adder_inst.intermediateResult2 ;
  wire \adder[3].adder_inst.intermediateResult3 ;
  wire \adder[3].adder_inst.out_carry ;
  wire \adder[3].adder_inst.out_sum ;
  wire \adder[4].adder_inst.in_A ;
  wire \adder[4].adder_inst.in_B ;
  wire \adder[4].adder_inst.in_carry ;
  wire \adder[4].adder_inst.intermediateResult1 ;
  wire \adder[4].adder_inst.intermediateResult2 ;
  wire \adder[4].adder_inst.intermediateResult3 ;
  wire \adder[4].adder_inst.out_carry ;
  wire \adder[4].adder_inst.out_sum ;
  wire \adder[5].adder_inst.in_A ;
  wire \adder[5].adder_inst.in_B ;
  wire \adder[5].adder_inst.in_carry ;
  wire \adder[5].adder_inst.intermediateResult1 ;
  wire \adder[5].adder_inst.intermediateResult2 ;
  wire \adder[5].adder_inst.intermediateResult3 ;
  wire \adder[5].adder_inst.out_carry ;
  wire \adder[5].adder_inst.out_sum ;
  wire \adder[6].adder_inst.in_A ;
  wire \adder[6].adder_inst.in_B ;
  wire \adder[6].adder_inst.in_carry ;
  wire \adder[6].adder_inst.intermediateResult1 ;
  wire \adder[6].adder_inst.intermediateResult2 ;
  wire \adder[6].adder_inst.intermediateResult3 ;
  wire \adder[6].adder_inst.out_carry ;
  wire \adder[6].adder_inst.out_sum ;
  wire \adder[7].adder_inst.in_A ;
  wire \adder[7].adder_inst.in_B ;
  wire \adder[7].adder_inst.in_carry ;
  wire \adder[7].adder_inst.intermediateResult1 ;
  wire \adder[7].adder_inst.intermediateResult2 ;
  wire \adder[7].adder_inst.intermediateResult3 ;
  wire \adder[7].adder_inst.out_carry ;
  wire \adder[7].adder_inst.out_sum ;
  wire \adder[8].adder_inst.in_A ;
  wire \adder[8].adder_inst.in_B ;
  wire \adder[8].adder_inst.in_carry ;
  wire \adder[8].adder_inst.intermediateResult1 ;
  wire \adder[8].adder_inst.intermediateResult2 ;
  wire \adder[8].adder_inst.intermediateResult3 ;
  wire \adder[8].adder_inst.out_carry ;
  wire \adder[8].adder_inst.out_sum ;
  wire \adder[9].adder_inst.in_A ;
  wire \adder[9].adder_inst.in_B ;
  wire \adder[9].adder_inst.in_carry ;
  wire \adder[9].adder_inst.intermediateResult1 ;
  wire \adder[9].adder_inst.intermediateResult2 ;
  wire \adder[9].adder_inst.intermediateResult3 ;
  wire \adder[9].adder_inst.out_carry ;
  wire \adder[9].adder_inst.out_sum ;
  wire \carry[0] ;
  wire \carry[10] ;
  wire \carry[11] ;
  wire \carry[12] ;
  wire \carry[13] ;
  wire \carry[14] ;
  wire \carry[15] ;
  wire \carry[16] ;
  wire \carry[17] ;
  wire \carry[18] ;
  wire \carry[19] ;
  wire \carry[1] ;
  wire \carry[20] ;
  wire \carry[21] ;
  wire \carry[22] ;
  wire \carry[23] ;
  wire \carry[24] ;
  wire \carry[25] ;
  wire \carry[26] ;
  wire \carry[27] ;
  wire \carry[28] ;
  wire \carry[29] ;
  wire \carry[2] ;
  wire \carry[30] ;
  wire \carry[31] ;
  wire \carry[32] ;
  wire \carry[3] ;
  wire \carry[4] ;
  wire \carry[5] ;
  wire \carry[6] ;
  wire \carry[7] ;
  wire \carry[8] ;
  wire \carry[9] ;
  input [31:0] input_A;
  input [31:0] input_B;
  output [32:0] output_sum;
  assign \adder[0].adder_inst.intermediateResult1  = input_A[0] ^ input_B[0];
  assign \adder[0].adder_inst.intermediateResult3  = input_A[0] & input_B[0];
  assign \adder[10].adder_inst.intermediateResult1  = input_A[10] ^ input_B[10];
  assign \adder[10].adder_inst.intermediateResult2  = \adder[10].adder_inst.intermediateResult1  & \adder[10].adder_inst.in_carry ;
  assign \adder[10].adder_inst.intermediateResult3  = input_A[10] & input_B[10];
  assign \adder[10].adder_inst.out_sum  = \adder[10].adder_inst.intermediateResult1  ^ \adder[10].adder_inst.in_carry ;
  assign \adder[10].adder_inst.out_carry  = \adder[10].adder_inst.intermediateResult2  | \adder[10].adder_inst.intermediateResult3 ;
  assign \adder[11].adder_inst.intermediateResult1  = input_A[11] ^ input_B[11];
  assign \adder[11].adder_inst.intermediateResult2  = \adder[11].adder_inst.intermediateResult1  & \adder[10].adder_inst.out_carry ;
  assign \adder[11].adder_inst.intermediateResult3  = input_A[11] & input_B[11];
  assign \adder[11].adder_inst.out_sum  = \adder[11].adder_inst.intermediateResult1  ^ \adder[10].adder_inst.out_carry ;
  assign \adder[11].adder_inst.out_carry  = \adder[11].adder_inst.intermediateResult2  | \adder[11].adder_inst.intermediateResult3 ;
  assign \adder[12].adder_inst.intermediateResult1  = input_A[12] ^ input_B[12];
  assign \adder[12].adder_inst.intermediateResult2  = \adder[12].adder_inst.intermediateResult1  & \adder[11].adder_inst.out_carry ;
  assign \adder[12].adder_inst.intermediateResult3  = input_A[12] & input_B[12];
  assign \adder[12].adder_inst.out_sum  = \adder[12].adder_inst.intermediateResult1  ^ \adder[11].adder_inst.out_carry ;
  assign \adder[12].adder_inst.out_carry  = \adder[12].adder_inst.intermediateResult2  | \adder[12].adder_inst.intermediateResult3 ;
  assign \adder[13].adder_inst.intermediateResult1  = input_A[13] ^ input_B[13];
  assign \adder[13].adder_inst.intermediateResult2  = \adder[13].adder_inst.intermediateResult1  & \adder[12].adder_inst.out_carry ;
  assign \adder[13].adder_inst.intermediateResult3  = input_A[13] & input_B[13];
  assign \adder[13].adder_inst.out_sum  = \adder[13].adder_inst.intermediateResult1  ^ \adder[12].adder_inst.out_carry ;
  assign \adder[13].adder_inst.out_carry  = \adder[13].adder_inst.intermediateResult2  | \adder[13].adder_inst.intermediateResult3 ;
  assign \adder[14].adder_inst.intermediateResult1  = input_A[14] ^ input_B[14];
  assign \adder[14].adder_inst.intermediateResult2  = \adder[14].adder_inst.intermediateResult1  & \adder[13].adder_inst.out_carry ;
  assign \adder[14].adder_inst.intermediateResult3  = input_A[14] & input_B[14];
  assign \adder[14].adder_inst.out_sum  = \adder[14].adder_inst.intermediateResult1  ^ \adder[13].adder_inst.out_carry ;
  assign \adder[14].adder_inst.out_carry  = \adder[14].adder_inst.intermediateResult2  | \adder[14].adder_inst.intermediateResult3 ;
  assign \adder[15].adder_inst.intermediateResult1  = input_A[15] ^ input_B[15];
  assign \adder[15].adder_inst.intermediateResult2  = \adder[15].adder_inst.intermediateResult1  & \adder[14].adder_inst.out_carry ;
  assign \adder[15].adder_inst.intermediateResult3  = input_A[15] & input_B[15];
  assign \adder[15].adder_inst.out_sum  = \adder[15].adder_inst.intermediateResult1  ^ \adder[14].adder_inst.out_carry ;
  assign \adder[15].adder_inst.out_carry  = \adder[15].adder_inst.intermediateResult2  | \adder[15].adder_inst.intermediateResult3 ;
  assign \adder[16].adder_inst.intermediateResult1  = input_A[16] ^ input_B[16];
  assign \adder[16].adder_inst.intermediateResult2  = \adder[16].adder_inst.intermediateResult1  & \adder[15].adder_inst.out_carry ;
  assign \adder[16].adder_inst.intermediateResult3  = input_A[16] & input_B[16];
  assign \adder[16].adder_inst.out_sum  = \adder[16].adder_inst.intermediateResult1  ^ \adder[15].adder_inst.out_carry ;
  assign \adder[16].adder_inst.out_carry  = \adder[16].adder_inst.intermediateResult2  | \adder[16].adder_inst.intermediateResult3 ;
  assign \adder[17].adder_inst.intermediateResult1  = input_A[17] ^ input_B[17];
  assign \adder[17].adder_inst.intermediateResult2  = \adder[17].adder_inst.intermediateResult1  & \adder[16].adder_inst.out_carry ;
  assign \adder[17].adder_inst.intermediateResult3  = input_A[17] & input_B[17];
  assign \adder[17].adder_inst.out_sum  = \adder[17].adder_inst.intermediateResult1  ^ \adder[16].adder_inst.out_carry ;
  assign \adder[17].adder_inst.out_carry  = \adder[17].adder_inst.intermediateResult2  | \adder[17].adder_inst.intermediateResult3 ;
  assign \adder[18].adder_inst.intermediateResult1  = input_A[18] ^ input_B[18];
  assign \adder[18].adder_inst.intermediateResult2  = \adder[18].adder_inst.intermediateResult1  & \adder[17].adder_inst.out_carry ;
  assign \adder[18].adder_inst.intermediateResult3  = input_A[18] & input_B[18];
  assign \adder[18].adder_inst.out_sum  = \adder[18].adder_inst.intermediateResult1  ^ \adder[17].adder_inst.out_carry ;
  assign \adder[18].adder_inst.out_carry  = \adder[18].adder_inst.intermediateResult2  | \adder[18].adder_inst.intermediateResult3 ;
  assign \adder[19].adder_inst.intermediateResult1  = input_A[19] ^ input_B[19];
  assign \adder[19].adder_inst.intermediateResult2  = \adder[19].adder_inst.intermediateResult1  & \adder[18].adder_inst.out_carry ;
  assign \adder[19].adder_inst.intermediateResult3  = input_A[19] & input_B[19];
  assign \adder[19].adder_inst.out_sum  = \adder[19].adder_inst.intermediateResult1  ^ \adder[18].adder_inst.out_carry ;
  assign \adder[19].adder_inst.out_carry  = \adder[19].adder_inst.intermediateResult2  | \adder[19].adder_inst.intermediateResult3 ;
  assign \adder[1].adder_inst.intermediateResult1  = input_A[1] ^ input_B[1];
  assign \adder[1].adder_inst.intermediateResult2  = \adder[1].adder_inst.intermediateResult1  & \adder[0].adder_inst.intermediateResult3 ;
  assign \adder[1].adder_inst.intermediateResult3  = input_A[1] & input_B[1];
  assign \adder[1].adder_inst.out_sum  = \adder[1].adder_inst.intermediateResult1  ^ \adder[0].adder_inst.intermediateResult3 ;
  assign \adder[1].adder_inst.out_carry  = \adder[1].adder_inst.intermediateResult2  | \adder[1].adder_inst.intermediateResult3 ;
  assign \adder[20].adder_inst.intermediateResult1  = input_A[20] ^ input_B[20];
  assign \adder[20].adder_inst.intermediateResult2  = \adder[20].adder_inst.intermediateResult1  & \adder[19].adder_inst.out_carry ;
  assign \adder[20].adder_inst.intermediateResult3  = input_A[20] & input_B[20];
  assign \adder[20].adder_inst.out_sum  = \adder[20].adder_inst.intermediateResult1  ^ \adder[19].adder_inst.out_carry ;
  assign \adder[20].adder_inst.out_carry  = \adder[20].adder_inst.intermediateResult2  | \adder[20].adder_inst.intermediateResult3 ;
  assign \adder[21].adder_inst.intermediateResult1  = input_A[21] ^ input_B[21];
  assign \adder[21].adder_inst.intermediateResult2  = \adder[21].adder_inst.intermediateResult1  & \adder[20].adder_inst.out_carry ;
  assign \adder[21].adder_inst.intermediateResult3  = input_A[21] & input_B[21];
  assign \adder[21].adder_inst.out_sum  = \adder[21].adder_inst.intermediateResult1  ^ \adder[20].adder_inst.out_carry ;
  assign \adder[21].adder_inst.out_carry  = \adder[21].adder_inst.intermediateResult2  | \adder[21].adder_inst.intermediateResult3 ;
  assign \adder[22].adder_inst.intermediateResult1  = input_A[22] ^ input_B[22];
  assign \adder[22].adder_inst.intermediateResult2  = \adder[22].adder_inst.intermediateResult1  & \adder[21].adder_inst.out_carry ;
  assign \adder[22].adder_inst.intermediateResult3  = input_A[22] & input_B[22];
  assign \adder[22].adder_inst.out_sum  = \adder[22].adder_inst.intermediateResult1  ^ \adder[21].adder_inst.out_carry ;
  assign \adder[22].adder_inst.out_carry  = \adder[22].adder_inst.intermediateResult2  | \adder[22].adder_inst.intermediateResult3 ;
  assign \adder[23].adder_inst.intermediateResult1  = input_A[23] ^ input_B[23];
  assign \adder[23].adder_inst.intermediateResult2  = \adder[23].adder_inst.intermediateResult1  & \adder[22].adder_inst.out_carry ;
  assign \adder[23].adder_inst.intermediateResult3  = input_A[23] & input_B[23];
  assign \adder[23].adder_inst.out_sum  = \adder[23].adder_inst.intermediateResult1  ^ \adder[22].adder_inst.out_carry ;
  assign \adder[23].adder_inst.out_carry  = \adder[23].adder_inst.intermediateResult2  | \adder[23].adder_inst.intermediateResult3 ;
  assign \adder[24].adder_inst.intermediateResult1  = input_A[24] ^ input_B[24];
  assign \adder[24].adder_inst.intermediateResult2  = \adder[24].adder_inst.intermediateResult1  & \adder[23].adder_inst.out_carry ;
  assign \adder[24].adder_inst.intermediateResult3  = input_A[24] & input_B[24];
  assign \adder[24].adder_inst.out_sum  = \adder[24].adder_inst.intermediateResult1  ^ \adder[23].adder_inst.out_carry ;
  assign \adder[24].adder_inst.out_carry  = \adder[24].adder_inst.intermediateResult2  | \adder[24].adder_inst.intermediateResult3 ;
  assign \adder[25].adder_inst.intermediateResult1  = input_A[25] ^ input_B[25];
  assign \adder[25].adder_inst.intermediateResult2  = \adder[25].adder_inst.intermediateResult1  & \adder[24].adder_inst.out_carry ;
  assign \adder[25].adder_inst.intermediateResult3  = input_A[25] & input_B[25];
  assign \adder[25].adder_inst.out_sum  = \adder[25].adder_inst.intermediateResult1  ^ \adder[24].adder_inst.out_carry ;
  assign \adder[25].adder_inst.out_carry  = \adder[25].adder_inst.intermediateResult2  | \adder[25].adder_inst.intermediateResult3 ;
  assign \adder[26].adder_inst.intermediateResult1  = input_A[26] ^ input_B[26];
  assign \adder[26].adder_inst.intermediateResult2  = \adder[26].adder_inst.intermediateResult1  & \adder[25].adder_inst.out_carry ;
  assign \adder[26].adder_inst.intermediateResult3  = input_A[26] & input_B[26];
  assign \adder[26].adder_inst.out_sum  = \adder[26].adder_inst.intermediateResult1  ^ \adder[25].adder_inst.out_carry ;
  assign \adder[26].adder_inst.out_carry  = \adder[26].adder_inst.intermediateResult2  | \adder[26].adder_inst.intermediateResult3 ;
  assign \adder[27].adder_inst.intermediateResult1  = input_A[27] ^ input_B[27];
  assign \adder[27].adder_inst.intermediateResult2  = \adder[27].adder_inst.intermediateResult1  & \adder[26].adder_inst.out_carry ;
  assign \adder[27].adder_inst.intermediateResult3  = input_A[27] & input_B[27];
  assign \adder[27].adder_inst.out_sum  = \adder[27].adder_inst.intermediateResult1  ^ \adder[26].adder_inst.out_carry ;
  assign \adder[27].adder_inst.out_carry  = \adder[27].adder_inst.intermediateResult2  | \adder[27].adder_inst.intermediateResult3 ;
  assign \adder[28].adder_inst.intermediateResult1  = input_A[28] ^ input_B[28];
  assign \adder[28].adder_inst.intermediateResult2  = \adder[28].adder_inst.intermediateResult1  & \adder[27].adder_inst.out_carry ;
  assign \adder[28].adder_inst.intermediateResult3  = input_A[28] & input_B[28];
  assign \adder[28].adder_inst.out_sum  = \adder[28].adder_inst.intermediateResult1  ^ \adder[27].adder_inst.out_carry ;
  assign \adder[28].adder_inst.out_carry  = \adder[28].adder_inst.intermediateResult2  | \adder[28].adder_inst.intermediateResult3 ;
  assign \adder[29].adder_inst.intermediateResult1  = input_A[29] ^ input_B[29];
  assign \adder[29].adder_inst.intermediateResult2  = \adder[29].adder_inst.intermediateResult1  & \adder[28].adder_inst.out_carry ;
  assign \adder[29].adder_inst.intermediateResult3  = input_A[29] & input_B[29];
  assign \adder[29].adder_inst.out_sum  = \adder[29].adder_inst.intermediateResult1  ^ \adder[28].adder_inst.out_carry ;
  assign \adder[29].adder_inst.out_carry  = \adder[29].adder_inst.intermediateResult2  | \adder[29].adder_inst.intermediateResult3 ;
  assign \adder[2].adder_inst.intermediateResult1  = input_A[2] ^ input_B[2];
  assign \adder[2].adder_inst.intermediateResult2  = \adder[2].adder_inst.intermediateResult1  & \adder[1].adder_inst.out_carry ;
  assign \adder[2].adder_inst.intermediateResult3  = input_A[2] & input_B[2];
  assign \adder[2].adder_inst.out_sum  = \adder[2].adder_inst.intermediateResult1  ^ \adder[1].adder_inst.out_carry ;
  assign \adder[2].adder_inst.out_carry  = \adder[2].adder_inst.intermediateResult2  | \adder[2].adder_inst.intermediateResult3 ;
  assign \adder[30].adder_inst.intermediateResult1  = input_A[30] ^ input_B[30];
  assign \adder[30].adder_inst.intermediateResult2  = \adder[30].adder_inst.intermediateResult1  & \adder[29].adder_inst.out_carry ;
  assign \adder[30].adder_inst.intermediateResult3  = input_A[30] & input_B[30];
  assign \adder[30].adder_inst.out_sum  = \adder[30].adder_inst.intermediateResult1  ^ \adder[29].adder_inst.out_carry ;
  assign \adder[30].adder_inst.out_carry  = \adder[30].adder_inst.intermediateResult2  | \adder[30].adder_inst.intermediateResult3 ;
  assign \adder[31].adder_inst.intermediateResult1  = input_A[31] ^ input_B[31];
  assign \adder[31].adder_inst.intermediateResult2  = \adder[31].adder_inst.intermediateResult1  & \adder[30].adder_inst.out_carry ;
  assign \adder[31].adder_inst.intermediateResult3  = input_A[31] & input_B[31];
  assign \adder[31].adder_inst.out_sum  = \adder[31].adder_inst.intermediateResult1  ^ \adder[30].adder_inst.out_carry ;
  assign \adder[31].adder_inst.out_carry  = \adder[31].adder_inst.intermediateResult2  | \adder[31].adder_inst.intermediateResult3 ;
  assign \adder[3].adder_inst.intermediateResult1  = input_A[3] ^ input_B[3];
  assign \adder[3].adder_inst.intermediateResult2  = \adder[3].adder_inst.intermediateResult1  & \adder[2].adder_inst.out_carry ;
  assign \adder[3].adder_inst.intermediateResult3  = input_A[3] & input_B[3];
  assign \adder[3].adder_inst.out_sum  = \adder[3].adder_inst.intermediateResult1  ^ \adder[2].adder_inst.out_carry ;
  assign \adder[3].adder_inst.out_carry  = \adder[3].adder_inst.intermediateResult2  | \adder[3].adder_inst.intermediateResult3 ;
  assign \adder[4].adder_inst.intermediateResult1  = input_A[4] ^ input_B[4];
  assign \adder[4].adder_inst.intermediateResult2  = \adder[4].adder_inst.intermediateResult1  & \adder[3].adder_inst.out_carry ;
  assign \adder[4].adder_inst.intermediateResult3  = input_A[4] & input_B[4];
  assign \adder[4].adder_inst.out_sum  = \adder[4].adder_inst.intermediateResult1  ^ \adder[3].adder_inst.out_carry ;
  assign \adder[4].adder_inst.out_carry  = \adder[4].adder_inst.intermediateResult2  | \adder[4].adder_inst.intermediateResult3 ;
  assign \adder[5].adder_inst.intermediateResult1  = input_A[5] ^ input_B[5];
  assign \adder[5].adder_inst.intermediateResult2  = \adder[5].adder_inst.intermediateResult1  & \adder[4].adder_inst.out_carry ;
  assign \adder[5].adder_inst.intermediateResult3  = input_A[5] & input_B[5];
  assign \adder[5].adder_inst.out_sum  = \adder[5].adder_inst.intermediateResult1  ^ \adder[4].adder_inst.out_carry ;
  assign \adder[5].adder_inst.out_carry  = \adder[5].adder_inst.intermediateResult2  | \adder[5].adder_inst.intermediateResult3 ;
  assign \adder[6].adder_inst.intermediateResult1  = input_A[6] ^ input_B[6];
  assign \adder[6].adder_inst.intermediateResult2  = \adder[6].adder_inst.intermediateResult1  & \adder[5].adder_inst.out_carry ;
  assign \adder[6].adder_inst.intermediateResult3  = input_A[6] & input_B[6];
  assign \adder[6].adder_inst.out_sum  = \adder[6].adder_inst.intermediateResult1  ^ \adder[5].adder_inst.out_carry ;
  assign \adder[6].adder_inst.out_carry  = \adder[6].adder_inst.intermediateResult2  | \adder[6].adder_inst.intermediateResult3 ;
  assign \adder[7].adder_inst.intermediateResult1  = input_A[7] ^ input_B[7];
  assign \adder[7].adder_inst.intermediateResult2  = \adder[7].adder_inst.intermediateResult1  & \adder[6].adder_inst.out_carry ;
  assign \adder[7].adder_inst.intermediateResult3  = input_A[7] & input_B[7];
  assign \adder[7].adder_inst.out_sum  = \adder[7].adder_inst.intermediateResult1  ^ \adder[6].adder_inst.out_carry ;
  assign \adder[7].adder_inst.out_carry  = \adder[7].adder_inst.intermediateResult2  | \adder[7].adder_inst.intermediateResult3 ;
  assign \adder[8].adder_inst.intermediateResult1  = input_A[8] ^ input_B[8];
  assign \adder[8].adder_inst.intermediateResult2  = \adder[8].adder_inst.intermediateResult1  & \adder[7].adder_inst.out_carry ;
  assign \adder[8].adder_inst.intermediateResult3  = input_A[8] & input_B[8];
  assign \adder[8].adder_inst.out_sum  = \adder[8].adder_inst.intermediateResult1  ^ \adder[7].adder_inst.out_carry ;
  assign \adder[8].adder_inst.out_carry  = \adder[8].adder_inst.intermediateResult2  | \adder[8].adder_inst.intermediateResult3 ;
  assign \adder[9].adder_inst.intermediateResult1  = input_A[9] ^ input_B[9];
  assign \adder[9].adder_inst.intermediateResult2  = \adder[9].adder_inst.intermediateResult1  & \adder[8].adder_inst.out_carry ;
  assign \adder[9].adder_inst.intermediateResult3  = input_A[9] & input_B[9];
  assign \adder[9].adder_inst.out_sum  = \adder[9].adder_inst.intermediateResult1  ^ \adder[8].adder_inst.out_carry ;
  assign \adder[10].adder_inst.in_carry  = \adder[9].adder_inst.intermediateResult2  | \adder[9].adder_inst.intermediateResult3 ;
  assign \adder[31].adder_inst.in_carry  = \adder[30].adder_inst.out_carry ;
  assign \adder[31].adder_inst.in_B  = input_B[31];
  assign \adder[31].adder_inst.in_A  = input_A[31];
  assign \adder[30].adder_inst.in_carry  = \adder[29].adder_inst.out_carry ;
  assign \adder[30].adder_inst.in_B  = input_B[30];
  assign \adder[30].adder_inst.in_A  = input_A[30];
  assign \adder[29].adder_inst.in_carry  = \adder[28].adder_inst.out_carry ;
  assign \adder[29].adder_inst.in_B  = input_B[29];
  assign \adder[29].adder_inst.in_A  = input_A[29];
  assign \adder[28].adder_inst.in_carry  = \adder[27].adder_inst.out_carry ;
  assign \adder[28].adder_inst.in_B  = input_B[28];
  assign \adder[28].adder_inst.in_A  = input_A[28];
  assign \adder[27].adder_inst.in_carry  = \adder[26].adder_inst.out_carry ;
  assign \adder[27].adder_inst.in_B  = input_B[27];
  assign \adder[27].adder_inst.in_A  = input_A[27];
  assign \adder[26].adder_inst.in_carry  = \adder[25].adder_inst.out_carry ;
  assign \adder[26].adder_inst.in_B  = input_B[26];
  assign \adder[26].adder_inst.in_A  = input_A[26];
  assign \adder[25].adder_inst.in_carry  = \adder[24].adder_inst.out_carry ;
  assign \adder[25].adder_inst.in_B  = input_B[25];
  assign \adder[25].adder_inst.in_A  = input_A[25];
  assign \adder[24].adder_inst.in_carry  = \adder[23].adder_inst.out_carry ;
  assign \adder[24].adder_inst.in_B  = input_B[24];
  assign \adder[24].adder_inst.in_A  = input_A[24];
  assign \adder[23].adder_inst.in_carry  = \adder[22].adder_inst.out_carry ;
  assign \adder[23].adder_inst.in_B  = input_B[23];
  assign \adder[23].adder_inst.in_A  = input_A[23];
  assign \adder[22].adder_inst.in_carry  = \adder[21].adder_inst.out_carry ;
  assign \adder[22].adder_inst.in_B  = input_B[22];
  assign \adder[22].adder_inst.in_A  = input_A[22];
  assign \adder[21].adder_inst.in_carry  = \adder[20].adder_inst.out_carry ;
  assign \adder[21].adder_inst.in_B  = input_B[21];
  assign \adder[21].adder_inst.in_A  = input_A[21];
  assign \adder[20].adder_inst.in_carry  = \adder[19].adder_inst.out_carry ;
  assign \adder[20].adder_inst.in_B  = input_B[20];
  assign \adder[20].adder_inst.in_A  = input_A[20];
  assign \adder[19].adder_inst.in_carry  = \adder[18].adder_inst.out_carry ;
  assign \adder[19].adder_inst.in_B  = input_B[19];
  assign \adder[19].adder_inst.in_A  = input_A[19];
  assign \adder[18].adder_inst.in_carry  = \adder[17].adder_inst.out_carry ;
  assign \adder[18].adder_inst.in_B  = input_B[18];
  assign \adder[18].adder_inst.in_A  = input_A[18];
  assign \adder[17].adder_inst.in_carry  = \adder[16].adder_inst.out_carry ;
  assign \adder[17].adder_inst.in_B  = input_B[17];
  assign \adder[17].adder_inst.in_A  = input_A[17];
  assign \adder[16].adder_inst.in_carry  = \adder[15].adder_inst.out_carry ;
  assign \adder[16].adder_inst.in_B  = input_B[16];
  assign \adder[16].adder_inst.in_A  = input_A[16];
  assign \adder[15].adder_inst.in_carry  = \adder[14].adder_inst.out_carry ;
  assign \adder[15].adder_inst.in_B  = input_B[15];
  assign \adder[15].adder_inst.in_A  = input_A[15];
  assign \adder[14].adder_inst.in_carry  = \adder[13].adder_inst.out_carry ;
  assign \adder[14].adder_inst.in_B  = input_B[14];
  assign \adder[14].adder_inst.in_A  = input_A[14];
  assign \adder[13].adder_inst.in_carry  = \adder[12].adder_inst.out_carry ;
  assign \adder[13].adder_inst.in_B  = input_B[13];
  assign \adder[13].adder_inst.in_A  = input_A[13];
  assign \adder[12].adder_inst.in_carry  = \adder[11].adder_inst.out_carry ;
  assign \adder[12].adder_inst.in_B  = input_B[12];
  assign \adder[12].adder_inst.in_A  = input_A[12];
  assign \adder[11].adder_inst.in_carry  = \adder[10].adder_inst.out_carry ;
  assign \adder[11].adder_inst.in_B  = input_B[11];
  assign \adder[11].adder_inst.in_A  = input_A[11];
  assign \adder[10].adder_inst.in_B  = input_B[10];
  assign \adder[10].adder_inst.in_A  = input_A[10];
  assign \adder[9].adder_inst.out_carry  = \adder[10].adder_inst.in_carry ;
  assign \adder[9].adder_inst.in_carry  = \adder[8].adder_inst.out_carry ;
  assign \adder[9].adder_inst.in_B  = input_B[9];
  assign \adder[9].adder_inst.in_A  = input_A[9];
  assign \adder[8].adder_inst.in_carry  = \adder[7].adder_inst.out_carry ;
  assign \adder[8].adder_inst.in_B  = input_B[8];
  assign \adder[8].adder_inst.in_A  = input_A[8];
  assign \adder[7].adder_inst.in_carry  = \adder[6].adder_inst.out_carry ;
  assign \adder[7].adder_inst.in_B  = input_B[7];
  assign \adder[7].adder_inst.in_A  = input_A[7];
  assign \adder[6].adder_inst.in_carry  = \adder[5].adder_inst.out_carry ;
  assign \adder[6].adder_inst.in_B  = input_B[6];
  assign \adder[6].adder_inst.in_A  = input_A[6];
  assign \adder[5].adder_inst.in_carry  = \adder[4].adder_inst.out_carry ;
  assign \adder[5].adder_inst.in_B  = input_B[5];
  assign \adder[5].adder_inst.in_A  = input_A[5];
  assign \adder[4].adder_inst.in_carry  = \adder[3].adder_inst.out_carry ;
  assign \adder[4].adder_inst.in_B  = input_B[4];
  assign \adder[4].adder_inst.in_A  = input_A[4];
  assign \adder[3].adder_inst.in_carry  = \adder[2].adder_inst.out_carry ;
  assign \adder[3].adder_inst.in_B  = input_B[3];
  assign \adder[3].adder_inst.in_A  = input_A[3];
  assign \adder[2].adder_inst.in_carry  = \adder[1].adder_inst.out_carry ;
  assign \adder[2].adder_inst.in_B  = input_B[2];
  assign \adder[2].adder_inst.in_A  = input_A[2];
  assign \adder[1].adder_inst.in_carry  = \adder[0].adder_inst.intermediateResult3 ;
  assign \adder[1].adder_inst.in_B  = input_B[1];
  assign \adder[1].adder_inst.in_A  = input_A[1];
  assign \adder[0].adder_inst.out_sum  = \adder[0].adder_inst.intermediateResult1 ;
  assign \adder[0].adder_inst.out_carry  = \adder[0].adder_inst.intermediateResult3 ;
  assign \adder[0].adder_inst.intermediateResult2  = 1'h0;
  assign \adder[0].adder_inst.in_carry  = 1'h0;
  assign \adder[0].adder_inst.in_B  = input_B[0];
  assign \adder[0].adder_inst.in_A  = input_A[0];
  assign \carry[0]  = 1'h0;
  assign \carry[10]  = \adder[10].adder_inst.in_carry ;
  assign \carry[11]  = \adder[10].adder_inst.out_carry ;
  assign \carry[12]  = \adder[11].adder_inst.out_carry ;
  assign \carry[13]  = \adder[12].adder_inst.out_carry ;
  assign \carry[14]  = \adder[13].adder_inst.out_carry ;
  assign \carry[15]  = \adder[14].adder_inst.out_carry ;
  assign \carry[16]  = \adder[15].adder_inst.out_carry ;
  assign \carry[17]  = \adder[16].adder_inst.out_carry ;
  assign \carry[18]  = \adder[17].adder_inst.out_carry ;
  assign \carry[19]  = \adder[18].adder_inst.out_carry ;
  assign \carry[1]  = \adder[0].adder_inst.intermediateResult3 ;
  assign \carry[20]  = \adder[19].adder_inst.out_carry ;
  assign \carry[21]  = \adder[20].adder_inst.out_carry ;
  assign \carry[22]  = \adder[21].adder_inst.out_carry ;
  assign \carry[23]  = \adder[22].adder_inst.out_carry ;
  assign \carry[24]  = \adder[23].adder_inst.out_carry ;
  assign \carry[25]  = \adder[24].adder_inst.out_carry ;
  assign \carry[26]  = \adder[25].adder_inst.out_carry ;
  assign \carry[27]  = \adder[26].adder_inst.out_carry ;
  assign \carry[28]  = \adder[27].adder_inst.out_carry ;
  assign \carry[29]  = \adder[28].adder_inst.out_carry ;
  assign \carry[2]  = \adder[1].adder_inst.out_carry ;
  assign \carry[30]  = \adder[29].adder_inst.out_carry ;
  assign \carry[31]  = \adder[30].adder_inst.out_carry ;
  assign \carry[32]  = \adder[31].adder_inst.out_carry ;
  assign \carry[3]  = \adder[2].adder_inst.out_carry ;
  assign \carry[4]  = \adder[3].adder_inst.out_carry ;
  assign \carry[5]  = \adder[4].adder_inst.out_carry ;
  assign \carry[6]  = \adder[5].adder_inst.out_carry ;
  assign \carry[7]  = \adder[6].adder_inst.out_carry ;
  assign \carry[8]  = \adder[7].adder_inst.out_carry ;
  assign \carry[9]  = \adder[8].adder_inst.out_carry ;
  assign output_sum = { \adder[31].adder_inst.out_carry , \adder[31].adder_inst.out_sum , \adder[30].adder_inst.out_sum , \adder[29].adder_inst.out_sum , \adder[28].adder_inst.out_sum , \adder[27].adder_inst.out_sum , \adder[26].adder_inst.out_sum , \adder[25].adder_inst.out_sum , \adder[24].adder_inst.out_sum , \adder[23].adder_inst.out_sum , \adder[22].adder_inst.out_sum , \adder[21].adder_inst.out_sum , \adder[20].adder_inst.out_sum , \adder[19].adder_inst.out_sum , \adder[18].adder_inst.out_sum , \adder[17].adder_inst.out_sum , \adder[16].adder_inst.out_sum , \adder[15].adder_inst.out_sum , \adder[14].adder_inst.out_sum , \adder[13].adder_inst.out_sum , \adder[12].adder_inst.out_sum , \adder[11].adder_inst.out_sum , \adder[10].adder_inst.out_sum , \adder[9].adder_inst.out_sum , \adder[8].adder_inst.out_sum , \adder[7].adder_inst.out_sum , \adder[6].adder_inst.out_sum , \adder[5].adder_inst.out_sum , \adder[4].adder_inst.out_sum , \adder[3].adder_inst.out_sum , \adder[2].adder_inst.out_sum , \adder[1].adder_inst.out_sum , \adder[0].adder_inst.intermediateResult1  };
endmodule
