module mhd_mit(a, b, f);
parameter _bit = 129;
parameter mhd = 48;
input [_bit - 1: 0] a;
input [_bit - 1: 0] b;
output f;
wire [_bit - 1: 0] diff;
wire [8: 0] sum;
assign diff[0] = a[0] ^ b[0];
assign diff[1] = a[1] ^ b[1];
assign diff[2] = a[2] ^ b[2];
assign diff[3] = a[3] ^ b[3];
assign diff[4] = a[4] ^ b[4];
assign diff[5] = a[5] ^ b[5];
assign diff[6] = a[6] ^ b[6];
assign diff[7] = a[7] ^ b[7];
assign diff[8] = a[8] ^ b[8];
assign diff[9] = a[9] ^ b[9];
assign diff[10] = a[10] ^ b[10];
assign diff[11] = a[11] ^ b[11];
assign diff[12] = a[12] ^ b[12];
assign diff[13] = a[13] ^ b[13];
assign diff[14] = a[14] ^ b[14];
assign diff[15] = a[15] ^ b[15];
assign diff[16] = a[16] ^ b[16];
assign diff[17] = a[17] ^ b[17];
assign diff[18] = a[18] ^ b[18];
assign diff[19] = a[19] ^ b[19];
assign diff[20] = a[20] ^ b[20];
assign diff[21] = a[21] ^ b[21];
assign diff[22] = a[22] ^ b[22];
assign diff[23] = a[23] ^ b[23];
assign diff[24] = a[24] ^ b[24];
assign diff[25] = a[25] ^ b[25];
assign diff[26] = a[26] ^ b[26];
assign diff[27] = a[27] ^ b[27];
assign diff[28] = a[28] ^ b[28];
assign diff[29] = a[29] ^ b[29];
assign diff[30] = a[30] ^ b[30];
assign diff[31] = a[31] ^ b[31];
assign diff[32] = a[32] ^ b[32];
assign diff[33] = a[33] ^ b[33];
assign diff[34] = a[34] ^ b[34];
assign diff[35] = a[35] ^ b[35];
assign diff[36] = a[36] ^ b[36];
assign diff[37] = a[37] ^ b[37];
assign diff[38] = a[38] ^ b[38];
assign diff[39] = a[39] ^ b[39];
assign diff[40] = a[40] ^ b[40];
assign diff[41] = a[41] ^ b[41];
assign diff[42] = a[42] ^ b[42];
assign diff[43] = a[43] ^ b[43];
assign diff[44] = a[44] ^ b[44];
assign diff[45] = a[45] ^ b[45];
assign diff[46] = a[46] ^ b[46];
assign diff[47] = a[47] ^ b[47];
assign diff[48] = a[48] ^ b[48];
assign diff[49] = a[49] ^ b[49];
assign diff[50] = a[50] ^ b[50];
assign diff[51] = a[51] ^ b[51];
assign diff[52] = a[52] ^ b[52];
assign diff[53] = a[53] ^ b[53];
assign diff[54] = a[54] ^ b[54];
assign diff[55] = a[55] ^ b[55];
assign diff[56] = a[56] ^ b[56];
assign diff[57] = a[57] ^ b[57];
assign diff[58] = a[58] ^ b[58];
assign diff[59] = a[59] ^ b[59];
assign diff[60] = a[60] ^ b[60];
assign diff[61] = a[61] ^ b[61];
assign diff[62] = a[62] ^ b[62];
assign diff[63] = a[63] ^ b[63];
assign diff[64] = a[64] ^ b[64];
assign diff[65] = a[65] ^ b[65];
assign diff[66] = a[66] ^ b[66];
assign diff[67] = a[67] ^ b[67];
assign diff[68] = a[68] ^ b[68];
assign diff[69] = a[69] ^ b[69];
assign diff[70] = a[70] ^ b[70];
assign diff[71] = a[71] ^ b[71];
assign diff[72] = a[72] ^ b[72];
assign diff[73] = a[73] ^ b[73];
assign diff[74] = a[74] ^ b[74];
assign diff[75] = a[75] ^ b[75];
assign diff[76] = a[76] ^ b[76];
assign diff[77] = a[77] ^ b[77];
assign diff[78] = a[78] ^ b[78];
assign diff[79] = a[79] ^ b[79];
assign diff[80] = a[80] ^ b[80];
assign diff[81] = a[81] ^ b[81];
assign diff[82] = a[82] ^ b[82];
assign diff[83] = a[83] ^ b[83];
assign diff[84] = a[84] ^ b[84];
assign diff[85] = a[85] ^ b[85];
assign diff[86] = a[86] ^ b[86];
assign diff[87] = a[87] ^ b[87];
assign diff[88] = a[88] ^ b[88];
assign diff[89] = a[89] ^ b[89];
assign diff[90] = a[90] ^ b[90];
assign diff[91] = a[91] ^ b[91];
assign diff[92] = a[92] ^ b[92];
assign diff[93] = a[93] ^ b[93];
assign diff[94] = a[94] ^ b[94];
assign diff[95] = a[95] ^ b[95];
assign diff[96] = a[96] ^ b[96];
assign diff[97] = a[97] ^ b[97];
assign diff[98] = a[98] ^ b[98];
assign diff[99] = a[99] ^ b[99];
assign diff[100] = a[100] ^ b[100];
assign diff[101] = a[101] ^ b[101];
assign diff[102] = a[102] ^ b[102];
assign diff[103] = a[103] ^ b[103];
assign diff[104] = a[104] ^ b[104];
assign diff[105] = a[105] ^ b[105];
assign diff[106] = a[106] ^ b[106];
assign diff[107] = a[107] ^ b[107];
assign diff[108] = a[108] ^ b[108];
assign diff[109] = a[109] ^ b[109];
assign diff[110] = a[110] ^ b[110];
assign diff[111] = a[111] ^ b[111];
assign diff[112] = a[112] ^ b[112];
assign diff[113] = a[113] ^ b[113];
assign diff[114] = a[114] ^ b[114];
assign diff[115] = a[115] ^ b[115];
assign diff[116] = a[116] ^ b[116];
assign diff[117] = a[117] ^ b[117];
assign diff[118] = a[118] ^ b[118];
assign diff[119] = a[119] ^ b[119];
assign diff[120] = a[120] ^ b[120];
assign diff[121] = a[121] ^ b[121];
assign diff[122] = a[122] ^ b[122];
assign diff[123] = a[123] ^ b[123];
assign diff[124] = a[124] ^ b[124];
assign diff[125] = a[125] ^ b[125];
assign diff[126] = a[126] ^ b[126];
assign diff[127] = a[127] ^ b[127];
assign diff[128] = a[128] ^ b[128];
assign sum = diff[0] + diff[1] + diff[2] + diff[3] + diff[4] + diff[5] + diff[6] + diff[7] + diff[8] + diff[9] + diff[10] + diff[11] + diff[12] + diff[13] + diff[14] + diff[15] + diff[16] + diff[17] + diff[18] + diff[19] + diff[20] + diff[21] + diff[22] + diff[23] + diff[24] + diff[25] + diff[26] + diff[27] + diff[28] + diff[29] + diff[30] + diff[31] + diff[32] + diff[33] + diff[34] + diff[35] + diff[36] + diff[37] + diff[38] + diff[39] + diff[40] + diff[41] + diff[42] + diff[43] + diff[44] + diff[45] + diff[46] + diff[47] + diff[48] + diff[49] + diff[50] + diff[51] + diff[52] + diff[53] + diff[54] + diff[55] + diff[56] + diff[57] + diff[58] + diff[59] + diff[60] + diff[61] + diff[62] + diff[63] + diff[64] + diff[65] + diff[66] + diff[67] + diff[68] + diff[69] + diff[70] + diff[71] + diff[72] + diff[73] + diff[74] + diff[75] + diff[76] + diff[77] + diff[78] + diff[79] + diff[80] + diff[81] + diff[82] + diff[83] + diff[84] + diff[85] + diff[86] + diff[87] + diff[88] + diff[89] + diff[90] + diff[91] + diff[92] + diff[93] + diff[94] + diff[95] + diff[96] + diff[97] + diff[98] + diff[99] + diff[100] + diff[101] + diff[102] + diff[103] + diff[104] + diff[105] + diff[106] + diff[107] + diff[108] + diff[109] + diff[110] + diff[111] + diff[112] + diff[113] + diff[114] + diff[115] + diff[116] + diff[117] + diff[118] + diff[119] + diff[120] + diff[121] + diff[122] + diff[123] + diff[124] + diff[125] + diff[126] + diff[127] + diff[128];
assign f = (sum > mhd);
endmodule
